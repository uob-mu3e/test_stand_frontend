-- megafunction wizard: %FIFO%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: dcfifo 

-- ============================================================
-- File Name: ip_dcfifo_mixed_widths.vhd
-- Megafunction Name(s):
--             dcfifo_mixed_widths
--
-- Simulation Library Files(s):
--             altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.0.0 Build 614 04/24/2018 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;


LIBRARY altera_mf;
USE altera_mf.all;

 
ENTITY ip_dcfifo_mixed_widths IS
    generic (
        ADDR_WIDTH_w    : positive := 8;
        DATA_WIDTH_w    : positive := 8;
        ADDR_WIDTH_r    : positive := 8;
        DATA_WIDTH_r    : positive := 8;
        SYNC_CLKS       : string := "TRUE";
        SHOWAHEAD       : string := "ON";
        REGOUT          : integer  := 1;
        DEVICE          : string := "Stratix IV"--;
    );
    PORT
    (
        aclr        : IN  STD_LOGIC  := '0';
        data        : IN  STD_LOGIC_VECTOR (DATA_WIDTH_w-1 DOWNTO 0);
        rdclk       : IN  STD_LOGIC;
        rdreq       : IN  STD_LOGIC;
        wrclk       : IN  STD_LOGIC;
        wrreq       : IN  STD_LOGIC;
        q           : OUT STD_LOGIC_VECTOR (DATA_WIDTH_r-1 DOWNTO 0);
        rdempty     : OUT STD_LOGIC;
        rdusedw     : OUT STD_LOGIC_VECTOR (ADDR_WIDTH_r-1 DOWNTO 0);
        wrfull      : OUT STD_LOGIC;
        wrusedw     : OUT STD_LOGIC_VECTOR (ADDR_WIDTH_w-1 DOWNTO 0)
    );
END ip_dcfifo_mixed_widths;


ARCHITECTURE SYN OF ip_dcfifo_mixed_widths IS

    SIGNAL sub_wire0    : STD_LOGIC_VECTOR (DATA_WIDTH_r-1 DOWNTO 0);
    SIGNAL sub_wire1    : STD_LOGIC;
    SIGNAL sub_wire2    : STD_LOGIC_VECTOR (ADDR_WIDTH_r-1 DOWNTO 0);
    SIGNAL sub_wire3    : STD_LOGIC;
    SIGNAL sub_wire4    : STD_LOGIC_VECTOR (ADDR_WIDTH_w-1 DOWNTO 0);

    COMPONENT dcfifo_mixed_widths
    GENERIC (
        clocks_are_synchronized    :   string;
        intended_device_family     :   string;
        lpm_numwords               :   natural;
        lpm_showahead              :   string;
        lpm_width                  :   natural;
        lpm_width_r                :   natural;
        lpm_widthu                 :   natural;
        lpm_widthu_r               :   natural;
        overflow_checking          :   string;
        rdsync_delaypipe           :   natural;
        read_aclr_synch            :   string;
        underflow_checking         :   string;
        use_eab                    :   string;
        write_aclr_synch           :   string;
        wrsync_delaypipe           :   natural--;
    );
    PORT (
        aclr        :   in  std_logic;
        data        :   in  std_logic_vector(DATA_WIDTH_w-1 downto 0);
        --eccstatus :   out std_logic_vector(2-1 downto 0);
        q           :   out std_logic_vector(DATA_WIDTH_r-1 downto 0);
        rdclk       :   in  std_logic;
        rdempty     :   out std_logic;
        --rdfull    :   out std_logic;
        rdreq       :   in  std_logic;
        rdusedw     :   out std_logic_vector(ADDR_WIDTH_r-1 downto 0);
        wrclk       :   in  std_logic;
        --wrempty   :   out std_logic;
        wrfull      :   out std_logic;
        wrreq       :   in  std_logic;
        wrusedw     :   out std_logic_vector(ADDR_WIDTH_w-1 downto 0)
    );
    END COMPONENT;

    signal rdusedw_reg : std_logic_vector(ADDR_WIDTH_r-1 downto 0);
    signal reset_n : std_logic;
    signal q0 : std_logic_vector(q'range);
    signal rdempty0 : std_logic;
    signal rdreq0, rdreq0_reg : std_logic;

BEGIN
    q0          <= sub_wire0(DATA_WIDTH_r-1 DOWNTO 0);
    rdempty0    <= sub_wire1;
    rdusedw     <= sub_wire2(ADDR_WIDTH_r-1 DOWNTO 0);

    process(rdclk, reset_n)
    begin
    if ( reset_n = '0' ) then
       rdusedw_reg  <= (others => '0');
       rdreq0_reg   <= '0';
    elsif ( rising_edge(rdclk) ) then
        rdusedw_reg <= rdusedw;
        rdreq0_reg <= rdreq0;
    end if;
    end process;

    wrfull      <= sub_wire3;
    wrusedw     <= sub_wire4(ADDR_WIDTH_w-1 DOWNTO 0);

    dcfifo_mixed_widths_component : dcfifo_mixed_widths
    GENERIC MAP (
        clocks_are_synchronized => SYNC_CLKS,
        intended_device_family  => DEVICE,
        lpm_numwords            => 2**ADDR_WIDTH_w,
        lpm_showahead           => SHOWAHEAD,
        lpm_width               => DATA_WIDTH_w,
        lpm_width_r             => DATA_WIDTH_r,
        lpm_widthu              => ADDR_WIDTH_w,
        lpm_widthu_r            => ADDR_WIDTH_r,
        overflow_checking       => "ON",
        rdsync_delaypipe        => 4,
        read_aclr_synch         => "ON",
        underflow_checking      => "ON",
        use_eab                 => "ON",
        write_aclr_synch        => "ON",
        wrsync_delaypipe        => 4
    )
    PORT MAP (
        aclr        => aclr,
        data        => data,
        rdclk       => rdclk,
        rdreq       => rdreq0,
        wrclk       => wrclk,
        wrreq       => wrreq,
        q           => sub_wire0,
        rdempty     => sub_wire1,
        rdusedw     => sub_wire2,
        wrfull      => sub_wire3,
        wrusedw     => sub_wire4
    );

    e_reset_n : entity work.reset_sync
    port map ( o_reset_n => reset_n, i_reset_n => not aclr, i_clk => rdclk );

    e_fifo_rreg : entity work.fifo_rreg
    generic map (
        g_N => work.util.value_if(SHOWAHEAD = "ON", REGOUT, 0),
        g_DATA_WIDTH => q'length--,
    )
    port map (
        o_rdata     => q,
        i_re        => rdreq,
        o_rempty    => rdempty,

        i_rdata     => q0,
        o_re        => rdreq0,
        i_rempty    => rdempty0,

        i_reset_n   => reset_n,
        i_clk       => rdclk--,
    );

END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
-- Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
-- Retrieval info: PRIVATE: AlmostFull NUMERIC "0"
-- Retrieval info: PRIVATE: AlmostFullThr NUMERIC "-1"
-- Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
-- Retrieval info: PRIVATE: Clock NUMERIC "4"
-- Retrieval info: PRIVATE: Depth NUMERIC "256"
-- Retrieval info: PRIVATE: Empty NUMERIC "1"
-- Retrieval info: PRIVATE: Full NUMERIC "1"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
-- Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
-- Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
-- Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
-- Retrieval info: PRIVATE: Optimize NUMERIC "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
-- Retrieval info: PRIVATE: UsedW NUMERIC "1"
-- Retrieval info: PRIVATE: Width NUMERIC "8"
-- Retrieval info: PRIVATE: dc_aclr NUMERIC "1"
-- Retrieval info: PRIVATE: diff_widths NUMERIC "0"
-- Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
-- Retrieval info: PRIVATE: output_width NUMERIC "8"
-- Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
-- Retrieval info: PRIVATE: rsFull NUMERIC "0"
-- Retrieval info: PRIVATE: rsUsedW NUMERIC "1"
-- Retrieval info: PRIVATE: sc_aclr NUMERIC "0"
-- Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
-- Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
-- Retrieval info: PRIVATE: wsFull NUMERIC "1"
-- Retrieval info: PRIVATE: wsUsedW NUMERIC "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "256"
-- Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "dcfifo"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "8"
-- Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
-- Retrieval info: CONSTANT: RDSYNC_DELAYPIPE NUMERIC "4"
-- Retrieval info: CONSTANT: READ_ACLR_SYNCH STRING "ON"
-- Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_ACLR_SYNCH STRING "ON"
-- Retrieval info: CONSTANT: WRSYNC_DELAYPIPE NUMERIC "4"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND "aclr"
-- Retrieval info: USED_PORT: data 0 0 8 0 INPUT NODEFVAL "data[7..0]"
-- Retrieval info: USED_PORT: q 0 0 8 0 OUTPUT NODEFVAL "q[7..0]"
-- Retrieval info: USED_PORT: rdclk 0 0 0 0 INPUT NODEFVAL "rdclk"
-- Retrieval info: USED_PORT: rdempty 0 0 0 0 OUTPUT NODEFVAL "rdempty"
-- Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL "rdreq"
-- Retrieval info: USED_PORT: rdusedw 0 0 8 0 OUTPUT NODEFVAL "rdusedw[7..0]"
-- Retrieval info: USED_PORT: wrclk 0 0 0 0 INPUT NODEFVAL "wrclk"
-- Retrieval info: USED_PORT: wrfull 0 0 0 0 OUTPUT NODEFVAL "wrfull"
-- Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL "wrreq"
-- Retrieval info: USED_PORT: wrusedw 0 0 8 0 OUTPUT NODEFVAL "wrusedw[7..0]"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: CONNECT: @data 0 0 8 0 data 0 0 8 0
-- Retrieval info: CONNECT: @rdclk 0 0 0 0 rdclk 0 0 0 0
-- Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
-- Retrieval info: CONNECT: @wrclk 0 0 0 0 wrclk 0 0 0 0
-- Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
-- Retrieval info: CONNECT: q 0 0 8 0 @q 0 0 8 0
-- Retrieval info: CONNECT: rdempty 0 0 0 0 @rdempty 0 0 0 0
-- Retrieval info: CONNECT: rdusedw 0 0 8 0 @rdusedw 0 0 8 0
-- Retrieval info: CONNECT: wrfull 0 0 0 0 @wrfull 0 0 0 0
-- Retrieval info: CONNECT: wrusedw 0 0 8 0 @wrusedw 0 0 8 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_dcfifo.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_dcfifo.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_dcfifo.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_dcfifo.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_dcfifo_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
