-- Sort hits by timestamp
-- New version for up to 45 input links and with memory for counter transmission
-- November 2019
-- niberger@uni-mainz.de

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;


use work.mupix.all;
use work.mudaq.all;

entity hitsorter_tb is
end hitsorter_tb;

architecture rtl of hitsorter_tb is

constant WRITECLK_PERIOD : time := 10 ns;
constant READCLK_PERIOD  : time := 8 ns;

signal		reset_n							: std_logic;										-- async reset
signal		writeclk						: std_logic;										-- clock for write/input side
signal 		tsclk							: std_logic;										-- clock for ts generation
signal		running							: std_logic;
signal		currentts						: ts_t;
signal		hit_in							: hit_array;
signal		hit_ena_in						: std_logic_vector(NCHIPS-1 downto 0);			-- valid hit
signal		readclk							: std_logic;										-- clock for read/output side
signal		data_out						: reg32;										-- packaged data out
signal		out_ena							: STD_LOGIC;									-- valid output data
signal		out_type						: std_logic_vector(3 downto 0);						
signal 		diagnostic_out					: sorter_reg_array;

begin


dut: entity work.hitsorter_wide 
	port map(
		reset_n							=> reset_n,
		writeclk						=> writeclk,
		running							=> running,
		currentts						=> currentts,
		hit_in							=> hit_in,
		hit_ena_in						=> hit_ena_in,
		readclk							=> readclk,
		data_out						=> data_out,
		out_ena							=> out_ena,
		out_type						=> out_type,
		diagnostic_out					=> diagnostic_out,
		delay							=> "01100000000"
		);

wclockgen: process
begin
	writeclk	<= '0';
	wait for WRITECLK_PERIOD/2;
	writeclk	<= '1';
	wait for WRITECLK_PERIOD/2;
end process;

tsclockgen: process
begin
	tsclk	<= '0';
	wait for WRITECLK_PERIOD/2;
	tsclk	<= '1';
	wait for WRITECLK_PERIOD/2;
end process;

rclockgen: process
begin
	readclk	<= '0';
	wait for READCLK_PERIOD/2;
	readclk	<= '1';
	wait for READCLK_PERIOD/2;
end process;

resetgen: process
begin
	reset_n <= '0';
	running <= '0';
	wait for 100 ns;
	reset_n	<= '1';
	wait for 100 ns;
	running <= '1';
	wait for 60000 ns;
	running <= '0';
	wait;
end process;

tsgen: process(reset_n, tsclk)
begin
if(reset_n = '0') then
	currentts	<= (others => '0');
elsif(tsclk'event and tsclk = '1') then
	if(running = '1') then
		currentts 	<= currentts + '1';
	end if;
end if;
end process;
	
hitgen: process
begin
	for i in NCHIPS-1 downto 0 loop
		hit_in(i)	<= (others => '0');
		hit_ena_in(i)	<= '0';
	end loop;
	wait for 30*WRITECLK_PERIOD;
	hit_in(0)		<= X"AAAAA001";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for 5*WRITECLK_PERIOD;
	hit_in(0)		<= X"BBBBB050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for 5*WRITECLK_PERIOD;
	hit_in(0)		<= X"CCCCC050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"DDDDD050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for 5*WRITECLK_PERIOD;
	hit_in(0)		<= X"EEEEE050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"11111050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for 5*WRITECLK_PERIOD;
	hit_in(0)		<= X"22222050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
	wait for 2*WRITECLK_PERIOD;
	hit_in(0)		<= X"33333050";
	hit_ena_in(0)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)		<= '0';
		
	wait for WRITECLK_PERIOD*100;
	hit_in(1)		<= X"BBBBB051";
	hit_ena_in(1)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"00000000";
	hit_ena_in(1)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(2)		<= X"CCCCC052";
	hit_ena_in(2)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(2)		<= X"00000000";
	hit_ena_in(2)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(3)		<= X"DDDDD053";
	hit_ena_in(3)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(3)		<= X"00000000";
	hit_ena_in(3)	<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(4)		<= X"EEEEE054";
	hit_ena_in(4)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(4)		<= X"00000000";
	hit_ena_in(4)	<= '0';
	wait for 5*WRITECLK_PERIOD;
	hit_in(5)		<= X"AAAAA055";
	hit_ena_in(5)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(5)		<= X"00000000";
	hit_ena_in(5)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(6)		<= X"BBBBB056";
	hit_ena_in(6)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(6)		<= X"00000000";
	hit_ena_in(6)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(7)		<= X"CCCCC057";
	hit_ena_in(7)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(7)		<= X"00000000";
	hit_ena_in(7)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(8)		<= X"DDDDD058";
	hit_ena_in(8)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(8)		<= X"00000000";
	hit_ena_in(8)	<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(9)		<= X"EEEEE059";
	hit_ena_in(9)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(9)		<= X"00000000";
	hit_ena_in(9)	<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(10)		<= X"BBBBB05A";
	hit_ena_in(10)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(10)		<= X"00000000";
	hit_ena_in(10)		<= '0';
	wait for WRITECLK_PERIOD;
	hit_in(11)		<= X"CCCCC05B";
	hit_ena_in(11)		<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(11)		<= X"00000000";
	hit_ena_in(11)		<= '0';
	wait for WRITECLK_PERIOD;
--	hit_in(12)		<= X"DDDDD07C";
--	hit_ena_in(12)		<= '1';
	wait for WRITECLK_PERIOD;
--	hit_in(12)		<= X"00000000";
--	hit_ena_in(12)	<= '0';
	wait for WRITECLK_PERIOD;
--	hit_in(13)		<= X"EEEEE07D";
--	hit_ena_in(13)		<= '1';
	wait for WRITECLK_PERIOD;
--	hit_in(13)		<= X"00000000";
--	hit_ena_in(13)	<= '0';
	wait for WRITECLK_PERIOD;
--	hit_in(14)		<= X"AAAAA07E";
--	hit_ena_in(14)		<= '1';
	wait for WRITECLK_PERIOD;
--	hit_in(14)		<= X"00000000";
--	hit_ena_in(14)	<= '0';
	wait for WRITECLK_PERIOD*5;
	hit_in(0)		<= X"00CCC080";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC080";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC080";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC080";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC080";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC080";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC080";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77BBB080";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC080";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC080";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC080";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC080";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC080";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC080";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC080";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	for i in 11 downto 0 loop
		hit_in(i)		<= X"00000000";
	end loop;
	hit_ena_in		<= (others => '0');
	wait for WRITECLK_PERIOD*5;
	hit_in(1)		<= X"11CCC085";
	hit_ena_in(1)	<= '1';
	hit_in(4)		<= X"44CCC085";
	hit_ena_in(4)	<= '1';
	hit_in(7)		<= X"77CCC085";
	hit_ena_in(7)	<= '1';
	hit_in(10)		<= X"aaCCC085";
	hit_ena_in(10)	<= '1';
--	hit_in(13)		<= X"ddCCC085";
--	hit_ena_in(13)	<= '1';
	wait for WRITECLK_PERIOD;
	for i in 11 downto 0 loop
		hit_in(i)		<= X"00000000";
	end loop;
	hit_ena_in		<= (others => '0');
	wait for WRITECLK_PERIOD*5;
	hit_in(0)		<= X"00DDD090";
	hit_ena_in(0)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00DDE090";
	hit_ena_in(0)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00DDF090";
	hit_ena_in(0)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in		<= (others => '0');
	wait for WRITECLK_PERIOD*5;
	hit_in(1)		<= X"11DD00BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD10BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD20BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD30BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD40BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD50BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD60BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD70BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD80BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DD90BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDA0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDB0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDC0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDD0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDE0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11DDF0BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"11EE10BF";
	hit_ena_in(1)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(1)		<= X"00000000";
	hit_ena_in		<= (others => '0');
	wait for WRITECLK_PERIOD*20;
	hit_in(0)		<= X"00CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77BBB180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"10CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"12CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"13CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"14CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"15CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"16CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"17CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"18CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"19CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"1aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"1bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"1cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"1dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"1eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"20CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"21CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"23CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"24CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"25CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"26CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"27CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"28CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"29CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"2aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"2bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"2cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"2dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"2eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"30CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"31CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"32CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"34CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"35CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"36CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"37CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"38CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"39CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"3aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"3bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"3cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"3dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"3eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"40CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"41CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"42CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"43CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"45CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"46CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"47CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"48CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"49CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"4aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"4bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"4cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"4dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"4eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"50CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"51CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"52CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"53CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"54CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"56CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"57CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"58CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"59CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"5aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"5bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"5cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"5dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"5eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"60CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"61CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"62CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"63CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"64CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"65CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"67CCC180";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"68CCC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"69CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"6aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"6bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"6cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"6dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"6eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC180";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"71CCC180";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"72CCC180";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"73CCC180";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"74CCC180";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"75CCC180";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"76CCC180";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CDC080";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"78CDC180";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"79CCC180";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"7aCCC180";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"7bCCC180";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"7cCCC180";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"7dCCC180";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"7eCCC180";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CDC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"10CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"12CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"13CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"14CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"15CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"16CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"17CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"18CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"19CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"1aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"1bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"1cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"1dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"1eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"20CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"21CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"23CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"24CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"25CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"26CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"27CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"28CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"29CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"2aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"2bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"2cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"2dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"2eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"30CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"31CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"32CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"34CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"35CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"36CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"37CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"38CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"39CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"3aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"3bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"3cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"3dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"3eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"40CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"41CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"42CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"43CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"45CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"46CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"47CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"48CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"49CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"4aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"4bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"4cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"4dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"4eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"50CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"51CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"52CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"53CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"54CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"56CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"57CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"58CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"59CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"5aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"5bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"5cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"5dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"5eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"60CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"61CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"62CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"63CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"64CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"65CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"67CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"68CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"69CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"6aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"6bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"6cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"6dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"6eCCC181";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC181";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"71CCC181";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"72CCC181";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"73CCC181";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"74CCC181";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"75CCC181";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"76CCC181";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CCC081";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"78CCC181";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"79CCC181";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"7aCCC181";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"7bCCC181";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"7cCCC181";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"7dCCC181";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"7eCCC181";
--	hit_ena_in(14)	<= '1';	
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CCC182";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"10CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"12CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"13CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"14CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"15CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"16CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"17CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"18CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"19CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"1aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"1bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"1cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"1dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"1eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"20CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"21CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"23CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"24CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"25CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"26CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"27CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"28CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"29CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"2aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"2bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"2cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"2dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"2eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"30CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"31CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"32CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"34CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"35CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"36CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"37CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"38CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"39CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"3aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"3bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"3cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"3dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"3eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"40CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"41CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"42CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"43CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"45CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"46CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"47CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"48CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"49CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"4aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"4bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"4cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"4dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"4eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"50CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"51CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"52CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"53CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"54CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"56CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"57CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"58CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"59CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"5aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"5bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"5cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"5dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"5eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"60CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"61CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"62CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"63CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"64CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"65CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"67CCC082";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"68CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"69CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"6aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"6bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"6cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"6dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"6eCCC182";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC182";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"71CCC182";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"72CCC182";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"73CCC182";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"74CCC182";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"75CCC182";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"76CCC182";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CBC182";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"78CCC182";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"79CCC182";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"7aCCC182";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"7bCCC182";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"7cCCC182";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"7dCCC182";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"7eCCC182";
--	hit_ena_in(14)	<= '1';	
		wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"10CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"12CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"13CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"14CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"15CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"16CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"17CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"18CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"19CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"1aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"1bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"1cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"1dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"1eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"20CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"21CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"23CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"24CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"25CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"26CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"27CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"28CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"29CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"2aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"2bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"2cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"2dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"2eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"30CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"31CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"32CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"34CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"35CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"36CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"37CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"38CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"39CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"3aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"3bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"3cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"3dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"3eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"40CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"41CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"42CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"43CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"45CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"46CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"47CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"48CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"49CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"4aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"4bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"4cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"4dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"4eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"50CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"51CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"52CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"53CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"54CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"56CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"57CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"58CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"59CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"5aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"5bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"5cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"5dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"5eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"60CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"61CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"62CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"63CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"64CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"65CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"67CCC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"68CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"69CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"6aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"6bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"6cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"6dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"6eCCC183";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC183";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"71CCC183";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"72CCC183";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"73CCC183";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"74CCC183";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"75CCC183";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"76CCC183";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CBC083";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"78CCC183";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"79CCC183";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"7aCCC183";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"7bCCC183";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"7cCCC183";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"7dCCC183";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"7eCCC183";
--	hit_ena_in(14)	<= '1';	
		wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"88CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"99CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"aaCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"bbCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"ccCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"ddCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"eeCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"10CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"11CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"12CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"13CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"14CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"15CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"16CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"17CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"18CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"19CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"1aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"1bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"1cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"1dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"1eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"20CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"21CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"22CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"23CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"24CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"25CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"26CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"27CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"28CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"29CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"2aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"2bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"2cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"2dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"2eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"30CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"31CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"32CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"33CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"34CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"35CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"36CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"37CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"38CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"39CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"3aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"3bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"3cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"3dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"3eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"40CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"41CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"42CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"43CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"44CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"45CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"46CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"47CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"48CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"49CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"4aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"4bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"4cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"4dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"4eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"50CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"51CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"52CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"53CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"54CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"55CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"56CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"57CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"58CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"59CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"5aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"5bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"5cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"5dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"5eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"60CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"61CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"62CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"63CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"64CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"65CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"66CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"67CCC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"68CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"69CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"6aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"6bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"6cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"6dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"6eCCC184";
--	hit_ena_in(14)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC184";
	hit_ena_in(0)	<= '1';
	hit_in(1)		<= X"71CCC184";
	hit_ena_in(1)	<= '1';
	hit_in(2)		<= X"72CCC184";
	hit_ena_in(2)	<= '1';
	hit_in(3)		<= X"73CCC184";
	hit_ena_in(3)	<= '1';
	hit_in(4)		<= X"74CCC184";
	hit_ena_in(4)	<= '1';
	hit_in(5)		<= X"75CCC184";
	hit_ena_in(5)	<= '1';
	hit_in(6)		<= X"76CCC184";
	hit_ena_in(6)	<= '1';
	hit_in(7)		<= X"77CBC084";
	hit_ena_in(7)	<= '1';
	hit_in(8)		<= X"78CCC184";
	hit_ena_in(8)	<= '1';
	hit_in(9)		<= X"79CCC184";
	hit_ena_in(9)	<= '1';
	hit_in(10)		<= X"7aCCC184";
	hit_ena_in(10)	<= '1';
	hit_in(11)		<= X"7bCCC184";
	hit_ena_in(11)	<= '1';
--	hit_in(12)		<= X"7cCCC184";
--	hit_ena_in(12)	<= '1';
--	hit_in(13)		<= X"7dCCC184";
--	hit_ena_in(13)	<= '1';
--	hit_in(14)		<= X"7eCCC184";
--	hit_ena_in(14)	<= '1';	
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"70CCC1A0";
	hit_ena_in(0)	<= '1';	
		wait for WRITECLK_PERIOD;
	for i in 11 downto 0 loop
		hit_in(i)		<= X"00000000";
	end loop;
	hit_ena_in		<= (others => '0');
    wait for 1900*WRITECLK_PERIOD;
	hit_in(0)		<= X"12345FFF";
	hit_ena_in(0)	<= '1';
	wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)	<= '0';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"ABAB0000";
	hit_ena_in(0)	<= '1';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)	<= '0';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"ABAB0007";
	hit_ena_in(0)	<= '1';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)	<= '0';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"ABAB0040";
	hit_ena_in(0)	<= '1';
    wait for WRITECLK_PERIOD;
	hit_in(0)		<= X"00000000";
	hit_ena_in(0)	<= '0';
	wait;
end process;

end architecture rtl;
