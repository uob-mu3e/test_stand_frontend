../a10_board/top.vhd