../../../fe_board/firmware/FEB_mutrig/lapse_counter.vhd