-- ip_madd.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
--library ip_madd_altera_fpdsp_block_180;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use ip_madd_altera_fpdsp_block_180.ip_madd_pkg.all;

entity ip_madd is
	port (
		aclr   : in  std_logic_vector(1 downto 0)  := (others => '0'); --   aclr.aclr
		ax     : in  std_logic_vector(31 downto 0) := (others => '0'); --     ax.ax
		ay     : in  std_logic_vector(31 downto 0) := (others => '0'); --     ay.ay
		az     : in  std_logic_vector(31 downto 0) := (others => '0'); --     az.az
		clk    : in  std_logic                     := '0';             --    clk.clk
		ena    : in  std_logic                     := '0';             --    ena.ena
		result : out std_logic_vector(31 downto 0)                     -- result.result
	);
end entity ip_madd;

architecture rtl of ip_madd is
begin

	fpdsp_block_0 : component work.ip_madd_altera_fpdsp_block_180_35ryh5a
		port map (
			clk    => clk,    --    clk.clk
			ena    => ena,    --    ena.ena
			aclr   => aclr,   --   aclr.aclr
			result => result, -- result.result
			ax     => ax,     --     ax.ax
			ay     => ay,     --     ay.ay
			az     => az      --     az.az
		);

end architecture rtl; -- of ip_madd
