../ddr3/ddr3_block.vhd