library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
entity f0_sim is
port(
data_feb0 : out std_logic_vector(31 downto 0);
datak_feb0 : out std_logic_vector(3 downto 0);
clk : in std_logic;
reset_n : in std_logic--;
);
end entity;
architecture behav of f0_sim is
begin
process
begin
if (reset_n = '0') then
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
else
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"000000bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"000d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c02e5382";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0eeb084";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"005fa284";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1ca3358";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0021f070";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"005f3810";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00656b70";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0042bffa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"004a3ea8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00ccb4c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"011eebfc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0164c000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01a30374";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01f799aa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0210fc7a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0259ad70";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"029726a4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02d4b60a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80261038";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80430234";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80683ee8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8058fcae";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80427eba";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80a0f8f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe46ee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"813b4ebc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8142e9e8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"819c5dec";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81c7107c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8201c758";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"826a7134";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8294ba86";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82c0be62";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f05e2106";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b147d2fa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1d02690";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b1597952";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"002c90d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00672590";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"006e1b20";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0040fdc4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0045facc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0081b83a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe084a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0109089a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"016f6752";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01b0f894";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01e52086";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02049820";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"025c5306";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02968ea0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02d0a63a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"801e8504";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80683ed8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"804f45c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8040fdc4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80478446";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80a715d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe474a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81095c84";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8152e088";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"818ae53e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81fd1f58";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"820cb898";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"825e53d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82a48648";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82c1fcd8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"4156d2d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"414752d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b14712c2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b15952d2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01777fd2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d15ed292";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f147c2c2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f06e27c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f06cfea0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f04db8a0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f07d7eb0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1e795a2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0001f37e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"007e7f94";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"004add48";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0042be2a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0041bd26";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00bb1afa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe706a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"011b6320";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0150296e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01affc5e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01dbe138";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"022ade9e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"026a3b60";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02a4a5ec";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02c888de";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"802a7be2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8047a974";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8043023e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80467bee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8042bfee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80b9f8f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe5888";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"810052fc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"816507c2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81a1877e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81ee3728";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"821ffeae";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8272dfac";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82a247ee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82cdc71a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70372aea";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70372aea";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"703b2aea";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f07a26e6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1c79160";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0005189a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"005f2410";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"006b26a0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00467dca";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0043bec4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00aaf9fc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe477c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0138353e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01556968";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01a3f3fa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01ccd084";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"023eb47c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"024f3760";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02b43946";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02c888fa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80311ef8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80430228";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8041ba4c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8049977e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8055ef7e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80be6fbc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe1fcc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8114b306";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"817cad28";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"818dd8a2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81e887ae";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8224eefc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82687e12";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"828d17c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82ee05ba";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2146d150";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a16912d0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"04e10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1c5f160";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00352b9e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"007dd7ba";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0058fca6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00423fe8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"005a0546";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0080b7c2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe57a0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"013a27a4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0175ed6c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"019f7ac6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01dcf724";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"020e7c7a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"027ab6c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02845afc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02d4b636";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80219a0a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8062d796";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8046b476";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"804bbb68";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80473734";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80ab9716";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe4d80";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8102cd6e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"816d6d2c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81ade1ee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81d85e28";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8222ef6e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82550a78";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82afc578";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82c1fcec";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0381fde";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1d757e2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0031c7f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00704200";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"004ef604";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0043fe9c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00467dde";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"008bbbb8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe70b2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"013d6ccc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"014ec1c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"018dfbbc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01cb27ca";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02103c3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"026a3b50";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02a0c0f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02c93b1c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"800efcfe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"805b1044";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80795b44";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80413f5a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80467bde";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8088f9f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80ccb4c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"811b168a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"814381c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81899c5c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81f8db8e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82353ef8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82706e5c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82ab2486";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82d4b62e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1f9e85e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"003692f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"007e7eba";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0047a976";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00507dbe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0041fef6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00bb5ab8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe1fe6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"011ab934";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01542d6e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01abf3c6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"01e287f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0233bdfc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"025ec43e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02850e50";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02c2b80a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0001";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"801e7df2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"804bd422";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"804f45d0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8043befc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8044fdbe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80af39f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80aeb8d8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80800000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe476c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"810b0284";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"815286a6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81b63598";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"81c839f0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8214c75c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"827dac24";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"828b01b4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"82c888ca";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0100";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"09620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0d620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe46f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe4744";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"11820000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"15820000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe46f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50fe0840";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"19a20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe475e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe58fe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"1dd10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80edc758";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe46f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b0fe4dbe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"21f10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"25f20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70fe4760";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2a010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe1f88";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0fe7004";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2e120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"36120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"40fe57fe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"90fe4772";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3a410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe583c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d0fe58dc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3e520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe4768";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"42720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50fe591c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0fe4ed8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"46a10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0fe70fc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d0fe08aa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70fe705e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"4ad20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe477e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50fe1f9c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"4ee20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"52e20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b0fe57de";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d0fe58f2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"57220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe4770";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"5b610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b0fe595c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"5f710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe468a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"63810000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe0850";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"67910000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe584e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe475e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"6be20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe593e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe1fe2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50fe082a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"90fe4d8c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe57ee";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d0fe58ea";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe475e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0fe085e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0ccb4c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"74720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"90fe70dc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"78920000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe4748";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20ccb4de";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7ca20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f125b9f6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"512b0a02";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80d10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe4756";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0edc74a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"85020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"60fe70be";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32067874";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"30ccb4dc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2397abe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"6210fc5c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21f2fac";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"89410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7231367e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2231be7e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70fe475a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f221bfbe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0fe5918";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21aba0a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"8d820000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe1f4c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe0874";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe1fa6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe4ef8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21f2fac";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f23dbe7e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"91f10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50f44074";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70fe4758";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0fe1fd2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe58b8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"96310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f03e478a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f03e4f8a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"703d3aac";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7038eaec";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a230be78";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"720e9c7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21f2fac";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3230b676";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62393e7e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a230a57e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"9aa20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b230b646";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe4744";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f1d757e2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e1c9840e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"421ac5c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c1c9c414";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"40fe57f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"9ed20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe4e82";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b219bc3e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe6fc0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"40fe5850";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3219bc0c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320ffc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21c80b4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320fc446";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f22cc480";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f23c4686";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"22017c7a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2207fc3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"221e0afa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"221e02fa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"223efc4a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320a5c3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"323082ca";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a3520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32308646";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7238a666";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"50fe469e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23384c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f23be4f4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"220ae060";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0fe1fcc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f2132fbc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8584";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"90fe7070";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2189084";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8086";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a7c20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"a0edd296";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e22118fc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"222632e4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f237f83e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62313a5a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62097c7a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"6201617a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62209a5a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21d38be";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2109090";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0866";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0fe4742";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2108686";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e0ccb4d8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe70d0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"ac510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f2132fbc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe7028";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21ac444";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe08bc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"30fe58e8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32289c76";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"322fbdfc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"72373a7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"921c4594";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"e20d7918";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0228d4b8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f23db4b8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21f2faa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"222e3cbc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3230b344";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"321e3b64";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"623ecc4c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3228b87c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b0b10000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"620ffc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7219bc3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b20ffc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"020bbc3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"021c4580";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3217fc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"723cfe3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320ffc7e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f20e2eae";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"123d61a4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b238b6f4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"021cc684";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3201647a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62209ae2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23b84d4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c80b4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d2019084";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3219bc3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe6fd6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b4e20000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe46f8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"322e7afa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe476e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"322e5afc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b9020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"80fe084c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21ac5c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21ac0c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8080";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"02108090";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3220d486";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"021cb580";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"221e3afa";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3219bc0a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"620a7c3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"0220d494";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23b84c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b20c80c4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b22cc484";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"023d8484";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe57dc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"bd620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23bc486";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe0876";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"40fe474c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"10fe4df2";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7219bc3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"2207fc0c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32017c7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"62107878";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"32263a7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b231bafc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2113a3a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b20db8b4";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8404";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f0fe57c8";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f221ba7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320ffc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3230be78";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"723bf800";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"d0ccb4d0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7219bc3e";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c2010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"020db086";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f21fd4de";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c6220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"20fe592c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"00fe4772";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8584";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b21c8584";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"020d8084";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"c0fe5f3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"620e7c7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"320f7c64";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"221a3c0c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"7238fe3c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"623b7abc";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f221ba7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"322f3e66";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23bc6b6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"722afdbe";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f22fb6e6";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"ca810000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"e8feb0bc";
datak_feb0 <= "0001";
wait until rising_edge(clk);
data_feb0 <= x"00000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"ce820000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc000000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc010000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc020000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc030000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc040000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc050000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc060000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc070000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc080000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc090000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc0f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc100000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"f03e478a";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc110000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc120000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc130000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc140000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc150000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc160000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc170000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc180000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc190000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc1f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc200000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc210000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc220000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc230000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc240000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc250000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc260000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc270000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc280000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc290000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"70382aec";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"3217fc7c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc2f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc300000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc310000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc320000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc330000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc340000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc350000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc360000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc370000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"321e843c";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc380000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc390000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc3f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc400000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc410000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc420000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc430000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc440000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc450000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc460000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc470000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc480000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc490000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc4f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc500000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc510000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc520000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc530000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc540000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc550000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc560000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc570000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc580000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc590000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc5f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc600000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc610000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc620000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc630000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc640000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc650000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc660000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc670000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc680000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc690000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc6f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc700000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc710000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc720000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc730000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc740000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc750000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc760000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc770000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc780000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b2108580";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"b23b84c0";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc790000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7a0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7b0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7c0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7d0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7e0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc7f0000";
datak_feb0 <= "0000";
wait until rising_edge(clk);
data_feb0 <= x"fc00009c";
datak_feb0 <= "0001";
wait until rising_edge(clk);
end if;
end process;
end architecture;
