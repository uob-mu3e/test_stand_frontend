../ddr3/ddr3_memory_controller.vhd