library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
entity f1_sim is
port(
data_feb1 : out std_logic_vector(31 downto 0);
datak_feb1 : out std_logic_vector(3 downto 0);
clk : in std_logic;
reset_n : in std_logic--;
);
end entity;
architecture behav of f1_sim is
begin
process
begin
if (reset_n = '0') then
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
else
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"000000bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"00100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"212da900";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e104320c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c00adc90";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0787272";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0e480f0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c10f6b08";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c11c79ec";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c14b6460";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c27bbd38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2b6c35c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c29dcf48";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2fb79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40086436";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4059773e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40e480fc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"411239b6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4119a79e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"416f66e6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"425d3c22";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42be4a0a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a80d0a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42e047e6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42b64a08";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a563a0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c03e08c6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c046c684";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c08f7d7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0e580ba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c101f902";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c104320c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c15dacdc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c18d242c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2773f8a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c29a8888";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c298e8f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2fb7e88";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"401e5420";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40780b4c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"408e7c42";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40e5808e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41173588";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"411821a6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41419434";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418eb8ae";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4247da9a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4297f090";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4292bcb8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42edff60";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a54ba0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c001fe04";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c065d3aa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0f98068";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1144cb0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c11332f6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1685c86";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1b31efe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2593c10";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2a4cb8a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c29f4acc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2edd8a2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4023d8c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"407bab62";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40e480c2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"410f3e38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"410b6f7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"417a769a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418dbd26";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"424a0402";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42ba2fde";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42828c0a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42e042c6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11dd6be";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ce94e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"04c10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c006a2ce";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c05c71c2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0990504";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0e58082";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c11d55ca";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1091a46";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c152c584";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c18e3c24";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2777c10";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2a33924";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2992a60";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2ecddba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40381520";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4044c1c8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40b043ac";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40bc4384";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40f80088";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4110c2bc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4105f57c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"414a7538";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418e3c24";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"426ead6c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a54b88";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42918c60";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42c10544";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c02626ea";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c06bb9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0f800ba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1143188";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1191ac2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c160490a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c26c080c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2b94584";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2a10924";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2eadf26";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"403691a2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"406ce82e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40bc7b9e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40e480e6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41128cca";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"411d1dbc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41614484";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418dac24";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42555286";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a0250c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a33be4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42e047c6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c04495d8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0e580b6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c118a386";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1067706";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c15a9d2c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c18e3c3c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c24d805e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2a9d522";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c296888c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2fd8dfe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"400c7ef4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40772f1e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40e58090";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"410e41c8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"411d6888";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41462184";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418be5bc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"424e1e1a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42b4150a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42a00e7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42d1e424";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c007afb0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0435fae";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c080bd78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c0f800aa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c11a51c2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1175dfa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1407cba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c18e2522";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c24e0246";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2ae0dd4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2890cbe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2fdb9f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4033f796";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"405338d6";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40af3bc2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40f800a2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4105b808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"410d2e06";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"414ab634";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"418e2522";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"41c00000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4266cf8e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42820a8e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42baeffe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"42d93e3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d1282740";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"09310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11dd6be";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ce94e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ebcc8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f113f7f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0d610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0f800b4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"111ff840";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"31214600";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d0f98058";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"70f6c0ce";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"11910000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11dd6be";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ce94e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ebcc8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f113f7f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"15d20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a12f06c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a13c2d80";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1220f40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e13c57c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"19e10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"1e110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"61313980";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"22210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"26510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0f8009a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"80d1c00c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b132f1c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"70e7001e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"2aa10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"90f80084";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"2ed20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"413b7bc0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"712d6a40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"70e480f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0d98972";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"90e58098";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"33120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"37220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b13867c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e12f43c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f130b8c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"3b610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0e580a2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"10d1c000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f251a164";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"326cb980";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"3fa20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"024d783c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f26a8c78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026af9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726af9a8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"72567c78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726bf9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24bbc3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"612b5240";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026afc38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25c3c3c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"027b79bc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"024c7c3c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"43f10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c26eb8b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0e480ec";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"90f9805a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"48310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d130f9c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f12a1b00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"4c420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7271f9fc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a25d2928";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"725a7c78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"724e7c78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7249d938";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"027b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"527b79a8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b4180";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726f39f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726f39f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79a8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"725c3c38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7262c9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"72583838";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b7990";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"027b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"126cf9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"126e469e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27b66a0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"50620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"3138d880";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"725c3c2c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27b79aa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"027b7998";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"54920000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f251a164";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a27e7938";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b120fac0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c1224e40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e12e6a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"58c10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0e480da";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a0d1c01e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"5d110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"513e2ac0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"613af9c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"612aa500";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"61120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"65420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0f8009a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"10e580b0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d1313940";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"69820000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"6db10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f251a164";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726f01f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b71b0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"2123b100";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"311e3f40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"413c3ac0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"713e1180";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"71e20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0e480ec";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"50f9c00e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e2448068";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27d26a4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"76320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0242b072";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"024d9baa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f251a164";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d7b82";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2487ffe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d7bba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d7e1a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d4382";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d7bba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b7988";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026af9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026cbc78";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b41b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7261f1f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"725f31f0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727b79b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726cf9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"72557bb8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a26e5b2a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27b66a0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27e6fae";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27e7f86";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"02527070";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a13898c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b1217a40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c133cdc0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"726cf9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"727c79bc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"725c3838";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25c3fbc";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026cf9b8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"72769bf8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7a720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026cfb92";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"827769ac";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"7ea10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c984a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"125bbbde";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"124e5e66";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"413aaf80";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"513d5680";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"512d6a40";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0e480da";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0d1c008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"82f20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"124e9e26";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"3259df5e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"87010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a1286200";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"8b110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f27d26a4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f26c2ba8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"926d427a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e26cbc1e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e26b9c5e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24e5fde";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24e1fde";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"8f710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25d3c3c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e25d3c38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131f808";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"93b10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11dd6be";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f252fd7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"026cdb9a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24c5fde";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e269da5e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"98010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2530c3c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f253b868";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f25f3838";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e26b9c5c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24c585c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24c585c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"824e1e5c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e26b9c62";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e275fb9c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c269dc58";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"9c620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c260a09e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e24d6626";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f251a164";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"525d1804";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a0a10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"21227a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1060a00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11dd6be";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ce94e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10ebcc8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f113f7f8";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1348b84";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a4f10000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1391980";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a9110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"713db848";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f26c212e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f2600386";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f26c292e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d25bbf10";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"325bbf3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"325bbf3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"325bbf3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f252fd7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"ad610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"324e5f7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"325bbf3e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"e2622c06";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"127e0f38";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"2122f000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"712be840";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f26d5c5c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b1a20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b5b20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"30f9c026";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"a13c7fc0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b139e1c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b120b940";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"b9d20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0b917fa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4544";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4544";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f09d3d04";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4544";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"be210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a043c4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c2310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f7d44";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f09d0524";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f09d0504";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"c6720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4542";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"408102c2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a07bc2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a043fa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a043c2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a043fa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1299900";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"cab20000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f10c2e7e";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f118a4fe";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11271f4";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f1113960";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"013dbc48";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"0131d008";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4544";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f09d0504";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f7d7c";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f7d44";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"d10e09e2";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"e8feb2bc";
datak_feb1 <= "0001";
wait until rising_edge(clk);
data_feb1 <= x"00000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"cf010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc000000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f0800000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc010000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f457a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4542";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f08f4542";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc020000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40a043fa";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc030000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc040000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc050000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc060000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc070000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc080000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc090000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc0f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc100000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc110000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc120000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc130000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc140000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc150000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc160000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc170000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc180000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc190000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"40ad43ba";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"f11f158a";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc1f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc200000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc210000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc220000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc230000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc240000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc250000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc260000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc270000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc280000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc290000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc2f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc300000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc310000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc320000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc330000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc340000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc350000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc360000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc370000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"51271f00";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"513432c0";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc380000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc390000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc3f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc400000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc410000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc420000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc430000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc440000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc450000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc460000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc470000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc480000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc490000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc4f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc500000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc510000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc520000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc530000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc540000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc550000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc560000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc570000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc580000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc590000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc5f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc600000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc610000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc620000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc630000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc640000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc650000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc660000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc670000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc680000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc690000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc6f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc700000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc710000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc720000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc730000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc740000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc750000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc760000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc770000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc780000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc790000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7a0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7b0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7c0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7d0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7e0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc7f0000";
datak_feb1 <= "0000";
wait until rising_edge(clk);
data_feb1 <= x"fc00009c";
datak_feb1 <= "0001";
wait until rising_edge(clk);
end if;
end process;
end architecture;
