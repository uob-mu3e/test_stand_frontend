library ieee;
use ieee.std_logic_1164.all;

package protocol is

    type data_merger_state is (idle, sending_data, sending_slowcontrol);
    --type feb_state is (idle, run_prep, sync, running, terminating, link_test, sync_test, reset_state, out_of_DAQ);

    constant HEADER_K:    std_logic_vector(31 downto 0) := x"000000bc";
    constant HEADER_K_DATAK:    std_logic_vector(3 downto 0) := "0001";
    constant WORD_ALIGN:    std_logic_vector(31 downto 0) := x"beefcafe";
    constant DATA_HEADER_ID:    std_logic_vector(5 downto 0) := "111010";
    constant DATA_SUB_HEADER_ID:    std_logic_vector(5 downto 0) := "111111";
    constant ACTIVE_SIGNAL_HEADER_ID:    std_logic_vector(5 downto 0) := "111101";
    constant RUN_TAIL_HEADER_ID:    std_logic_vector(5 downto 0) := "111110";
    constant TIMING_MEAS_HEADER_ID:    std_logic_vector(5 downto 0) := "111100";
    constant SC_HEADER_ID:    std_logic_vector(5 downto 0) := "111011";

end package protocol;

-- simple data generator (for slowcontrol and pixel data)
-- writes into pix_data_fifo and sc_data_fifo
-- only Header(sc or pix) + data
-- other headers/signals are added in data_merger.vhd

-- Martin Mueller, January 2019
-- Marius Koeppel, March 2019
-- Marius Koeppel, July 2019

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.protocol.all;


entity data_generator_a10_tb is
    port(
		clk:                 	in  std_logic;
		reset:               	in  std_logic;
		enable_pix:          	in  std_logic;
		random_seed:			in  std_logic_vector (15 downto 0);
		start_global_time:		in  std_logic_vector(47 downto 0);
		data_pix_generated:  	out std_logic_vector(31 downto 0);
		datak_pix_generated:  	out std_logic_vector(3 downto 0);
		data_pix_ready:      	out std_logic;
        slow_down:			    in  std_logic_vector(31 downto 0);
		state_out:  	        out std_logic_vector(3 downto 0)
);
end entity data_generator_a10_tb;

architecture rtl of data_generator_a10_tb is

component linear_shift is 
	generic (
		g_m             : integer           := 7;
		g_poly          : std_logic_vector  := "1100000" -- x^7+x^6+1 
	);
	port (
		i_clk           : in  std_logic;
		reset_n         : in  std_logic;
		i_sync_reset    : in  std_logic;
		i_seed          : in  std_logic_vector (g_m-1 downto 0);
		i_en            : in  std_logic;
		o_lsfr          : out std_logic_vector (g_m-1 downto 0)
	);
end component linear_shift;

----------------signals---------------------
	signal global_time:			  std_logic_vector(47 downto 0);
	signal reset_n:				  std_logic;
	-- state_types
	type data_header_states is (part1, part2, part3, part4, part5, trailer, overflow);
	signal data_header_state:   data_header_states;

	-- random signals
	signal lsfr_chip_id:     	  std_logic_vector (5 downto 0);
	signal lsfr_tot:     	  	  std_logic_vector (5 downto 0);
	signal lsfr_row:     	  	  std_logic_vector (7 downto 0);
	signal lsfr_col:     	     std_logic_vector (7 downto 0);
	signal lsfr_overflow:        std_logic_vector (15 downto 0);
	
	-- slow down signals
	signal waiting:				  std_logic;
	signal wait_counter:			  std_logic_vector(31 downto 0);

----------------begin data_generator------------------------
begin

	reset_n <= not reset;

	chip_id_shift : linear_shift
	generic map(
		g_m 	   		=> 6,
		g_poly 	   	=> "110000"
	)
	port map(
		i_clk    		=> clk,
		reset_n   		=> reset_n,
		i_sync_reset	=> reset,--sync_reset,
		i_seed   		=> random_seed(5 downto 0),
		i_en 				=> enable_pix,    
		o_lsfr 			=> lsfr_chip_id
	);
	
	pix_tot_shift : linear_shift
	generic map(
		g_m 	   		=> 6,
		g_poly 	   	=> "110000"
	)
	port map(
		i_clk    		=> clk,
		reset_n   		=> reset_n,
		i_sync_reset	=> reset,--sync_reset,
		i_seed   		=> random_seed(15 downto 10),
		i_en 				=> enable_pix,    
		o_lsfr 			=> lsfr_tot
	);
	
	pix_row_shift : linear_shift
	generic map(
		g_m 	   		=> 8,
		g_poly 	   	=> "10111000"
	)
	port map(
		i_clk    		=> clk,
		reset_n   		=> reset_n,
		i_sync_reset	=> reset,--sync_reset,
		i_seed   		=> random_seed(7 downto 0),
		i_en 				=> enable_pix,    
		o_lsfr 			=> lsfr_row
	);
	
	pix_col_shift : linear_shift
	generic map(
		g_m 	   		=> 8,
		g_poly 	   	=> "10111000"
	)
	port map(
		i_clk    		=> clk,
		reset_n   		=> reset_n,
		i_sync_reset	=> reset,--sync_reset,
		i_seed   		=> random_seed(8 downto 1),
		i_en 				=> enable_pix,    
		o_lsfr 			=> lsfr_col
	);
	
	overflow_shift : linear_shift
	generic map(
		g_m 	   		=> 16,
		g_poly 	   	=> "1101000000001000"
	)
	port map(
		i_clk    		=> clk,
		reset_n   		=> reset_n,
		i_sync_reset	=> reset,--sync_reset,
		i_seed   		=> random_seed,
		i_en 				=> enable_pix,    
		o_lsfr 			=> lsfr_overflow
	);

-- slow down process
process(clk, reset)
begin
	if(reset = '1' or enable_pix = '0') then
		waiting 			<= '0';
		wait_counter	<= (others => '0');
	elsif(rising_edge(clk)) then
		if(wait_counter >= slow_down) then
			wait_counter 	<= (others => '0');
			waiting 			<= '0';
		else
			wait_counter		<= wait_counter + '1';
			waiting			<= '1';
		end if;
	end if;
end process;
	
	
	
process (clk)

variable current_overflow : std_logic_vector(15 downto 0) := "0000000000000000";
variable overflow_idx	  : integer range 0 to 15 := 0;

begin
	if (reset = '1') then
		data_pix_ready          <= '0';
		--data_sc_ready           <= '0';
		data_pix_generated      <= (others => '0');
		--data_sc_generated       <= (others => '0');
		global_time       		<= start_global_time;
		--sc_data_counter         <= (others => '1');
		data_header_state			<= part1;
		--wait_cnt						<= (others => '0');
		current_overflow 			:= "0000000000000000";
		overflow_idx				:= 0;
	elsif rising_edge(clk) then
        -- generate pix data
        
        if(enable_pix = '1' and waiting = '0') then
				data_pix_ready <= '1';
				case data_header_state is
					when part1 =>
						state_out                         <= x"1";
						global_time                       <= global_time + '1';
						data_pix_generated(31 downto 26)  <= "111010";
						data_pix_generated(25 downto 8)   <= (others => '0');
						data_pix_generated(7 downto 0) 	  <= x"bc";
						datak_pix_generated               <= "0001";
						data_header_state 				  <= part2;
				
					when part2 =>
                        state_out <= x"2";
						data_pix_generated				    <= global_time(47 downto 16);
                        datak_pix_generated                 <= "0000";
						data_header_state 					<= part3;
					
					when part3 =>
						state_out <= x"3";
						data_pix_generated					<= global_time(15 downto 0) & x"0000";
						data_header_state 					<= part4;
						
					when part4 =>
						state_out <= x"4";
						data_pix_generated 					<= "0000" & DATA_SUB_HEADER_ID & global_time(9 downto 4) & lsfr_overflow;
						datak_pix_generated                 <= "0000";
						global_time							<= global_time + '1';
						overflow_idx 						:= 0;
						current_overflow					:= lsfr_overflow;
						data_header_state 					<= part5;
					
					when part5 =>
                        state_out <= x"5";
                        datak_pix_generated                 <= "0000";
						if (lsfr_chip_id = DATA_SUB_HEADER_ID) then
							data_pix_generated				<= "101010" & lsfr_row & lsfr_col & lsfr_tot;
						elsif (lsfr_chip_id = DATA_HEADER_ID) then
							data_pix_generated				<= "010101" & lsfr_row & lsfr_col & lsfr_tot;
						else
							data_pix_generated				<= lsfr_chip_id & lsfr_row & lsfr_col & lsfr_tot;
						end if;
						
						if (current_overflow(overflow_idx) = '1') then
							overflow_idx 						:= overflow_idx + 1;
							data_header_state					<= overflow;
						else
							overflow_idx 						:= overflow_idx + 1;
							global_time 						<= global_time + '1';
						end if;
						
						if (global_time(9 downto 0) = "1111111111") then
							data_header_state 				<= trailer;
						elsif (global_time(3 downto 0) = "1111") then
							data_header_state 				<= part4;
						end if;
							
					when overflow =>
						state_out <= x"6";
						datak_pix_generated                 <= "0000";
                        if (lsfr_chip_id = DATA_SUB_HEADER_ID) then
							data_pix_generated				<= "0000" & global_time(3 downto 0) & "000000" & global_time(21 downto 0);-- "101010" & lsfr_row & lsfr_col & lsfr_tot;
						elsif (lsfr_chip_id = DATA_HEADER_ID) then
							data_pix_generated				<= "0000" & global_time(3 downto 0) & "000000" & global_time(21 downto 0); -- "010101" & lsfr_row & lsfr_col & lsfr_tot;
						else
							data_pix_generated				<= "0000" & global_time(3 downto 0) & "000000" & global_time(21 downto 0); --lsfr_chip_id & lsfr_row & lsfr_col & lsfr_tot;
						end if;
						global_time 							<= global_time + '1';
						data_header_state						<= part5;
					
					when trailer =>
						state_out <= x"7";
						global_time <= global_time + '1';
						datak_pix_generated                 <= "0001";
						data_pix_generated(31 downto 8)	<= (others => '0');
						data_pix_generated(7 downto 0)	<= x"9c";
						data_header_state 					<= part1;
						
					when others =>
						state_out <= x"8";
						data_header_state 					<= trailer;
						---
				end case;
		else
			state_out <= x"F";
			data_pix_ready <= '0';
		end if;
    end if;
end process;



END rtl;
