----------------------------------------------------------------------------
-- storage for Mupix TDACs
-- M. Mueller, Feb 2022
-----------------------------------------------------------------------------

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

entity convert_col_row_reverse is
    port(
        i_addr  : in  std_logic_vector(8 downto 0);
        o_addr  : out std_logic_vector(8 downto 0)--;
    );
end entity convert_col_row_reverse;

architecture RTL of convert_col_row_reverse is

    signal mem_addr : std_logic_vector(11 downto 0);
    signal addr     : std_logic_vector(11 downto 0);

begin
    o_addr <= mem_addr(8 downto 0);
    addr   <= "000" & i_addr;

    process (addr) is
    begin
        case addr is  
            when x"135" => mem_addr <= x"00b";
            when x"0fa" => mem_addr <= x"00c";
            when x"136" => mem_addr <= x"00d";
            when x"0fb" => mem_addr <= x"00e";
            when x"137" => mem_addr <= x"00f";
            when x"0fc" => mem_addr <= x"010";
            when x"138" => mem_addr <= x"011";
            when x"0fd" => mem_addr <= x"012";
            when x"139" => mem_addr <= x"013";
            when x"0fe" => mem_addr <= x"014";
            when x"13a" => mem_addr <= x"015";
            when x"0ff" => mem_addr <= x"016";
            when x"13b" => mem_addr <= x"017";
            when x"100" => mem_addr <= x"018";
            when x"13c" => mem_addr <= x"019";
            when x"101" => mem_addr <= x"01a";
            when x"13d" => mem_addr <= x"01b";
            when x"102" => mem_addr <= x"01c";
            when x"13e" => mem_addr <= x"01d";
            when x"103" => mem_addr <= x"01e";
            when x"13f" => mem_addr <= x"01f";
            when x"104" => mem_addr <= x"020";
            when x"140" => mem_addr <= x"021";
            when x"105" => mem_addr <= x"022";
            when x"141" => mem_addr <= x"023";
            when x"106" => mem_addr <= x"024";
            when x"142" => mem_addr <= x"025";
            when x"107" => mem_addr <= x"026";
            when x"143" => mem_addr <= x"027";
            when x"108" => mem_addr <= x"028";
            when x"144" => mem_addr <= x"029";
            when x"109" => mem_addr <= x"02a";
            when x"145" => mem_addr <= x"02b";
            when x"10a" => mem_addr <= x"02c";
            when x"146" => mem_addr <= x"02d";
            when x"10b" => mem_addr <= x"02e";
            when x"147" => mem_addr <= x"02f";
            when x"10c" => mem_addr <= x"030";
            when x"148" => mem_addr <= x"031";
            when x"10d" => mem_addr <= x"032";
            when x"149" => mem_addr <= x"033";
            when x"10e" => mem_addr <= x"034";
            when x"14a" => mem_addr <= x"035";
            when x"10f" => mem_addr <= x"036";
            when x"14b" => mem_addr <= x"037";
            when x"110" => mem_addr <= x"038";
            when x"14c" => mem_addr <= x"039";
            when x"111" => mem_addr <= x"03a";
            when x"14d" => mem_addr <= x"03b";
            when x"112" => mem_addr <= x"03c";
            when x"14e" => mem_addr <= x"03d";
            when x"113" => mem_addr <= x"03e";
            when x"14f" => mem_addr <= x"03f";
            when x"114" => mem_addr <= x"040";
            when x"150" => mem_addr <= x"041";
            when x"115" => mem_addr <= x"042";
            when x"151" => mem_addr <= x"043";
            when x"116" => mem_addr <= x"044";
            when x"152" => mem_addr <= x"045";
            when x"117" => mem_addr <= x"046";
            when x"153" => mem_addr <= x"047";
            when x"118" => mem_addr <= x"048";
            when x"154" => mem_addr <= x"049";
            when x"119" => mem_addr <= x"04a";
            when x"155" => mem_addr <= x"04b";
            when x"11a" => mem_addr <= x"04c";
            when x"156" => mem_addr <= x"04d";
            when x"11b" => mem_addr <= x"04e";
            when x"157" => mem_addr <= x"04f";
            when x"11c" => mem_addr <= x"050";
            when x"158" => mem_addr <= x"051";
            when x"11d" => mem_addr <= x"052";
            when x"159" => mem_addr <= x"053";
            when x"11e" => mem_addr <= x"054";
            when x"15a" => mem_addr <= x"055";
            when x"11f" => mem_addr <= x"056";
            when x"15b" => mem_addr <= x"057";
            when x"120" => mem_addr <= x"058";
            when x"15c" => mem_addr <= x"059";
            when x"121" => mem_addr <= x"05a";
            when x"15d" => mem_addr <= x"05b";
            when x"122" => mem_addr <= x"05c";
            when x"15e" => mem_addr <= x"05d";
            when x"123" => mem_addr <= x"05e";
            when x"15f" => mem_addr <= x"05f";
            when x"124" => mem_addr <= x"060";
            when x"160" => mem_addr <= x"061";
            when x"125" => mem_addr <= x"062";
            when x"161" => mem_addr <= x"063";
            when x"126" => mem_addr <= x"064";
            when x"162" => mem_addr <= x"065";
            when x"127" => mem_addr <= x"066";
            when x"163" => mem_addr <= x"067";
            when x"128" => mem_addr <= x"068";
            when x"164" => mem_addr <= x"069";
            when x"129" => mem_addr <= x"06a";
            when x"165" => mem_addr <= x"06b";
            when x"12a" => mem_addr <= x"06c";
            when x"166" => mem_addr <= x"06d";
            when x"12b" => mem_addr <= x"06e";
            when x"167" => mem_addr <= x"06f";
            when x"12c" => mem_addr <= x"070";
            when x"168" => mem_addr <= x"071";
            when x"12d" => mem_addr <= x"072";
            when x"169" => mem_addr <= x"073";
            when x"12e" => mem_addr <= x"074";
            when x"16a" => mem_addr <= x"075";
            when x"12f" => mem_addr <= x"076";
            when x"16b" => mem_addr <= x"077";
            when x"130" => mem_addr <= x"078";
            when x"16c" => mem_addr <= x"079";
            when x"131" => mem_addr <= x"07a";
            when x"16d" => mem_addr <= x"07b";
            when x"132" => mem_addr <= x"07c";
            when x"16e" => mem_addr <= x"07d";
            when x"133" => mem_addr <= x"07e";
            when x"16f" => mem_addr <= x"07f";
            when x"134" => mem_addr <= x"080";
            when x"170" => mem_addr <= x"081";
            --when x"135" => mem_addr <= x"082"; -- Why does this show up again ?
            when x"03e" => mem_addr <= x"083";
            when x"000" => mem_addr <= x"084";
            when x"03f" => mem_addr <= x"085";
            when x"001" => mem_addr <= x"086";
            when x"040" => mem_addr <= x"087";
            when x"002" => mem_addr <= x"088";
            when x"041" => mem_addr <= x"089";
            when x"003" => mem_addr <= x"08a";
            when x"042" => mem_addr <= x"08b";
            when x"004" => mem_addr <= x"08c";
            when x"043" => mem_addr <= x"08d";
            when x"005" => mem_addr <= x"08e";
            when x"044" => mem_addr <= x"08f";
            when x"006" => mem_addr <= x"090";
            when x"045" => mem_addr <= x"091";
            when x"007" => mem_addr <= x"092";
            when x"046" => mem_addr <= x"093";
            when x"008" => mem_addr <= x"094";
            when x"047" => mem_addr <= x"095";
            when x"009" => mem_addr <= x"096";
            when x"048" => mem_addr <= x"097";
            when x"00a" => mem_addr <= x"098";
            when x"049" => mem_addr <= x"099";
            when x"00b" => mem_addr <= x"09a";
            when x"04a" => mem_addr <= x"09b";
            when x"00c" => mem_addr <= x"09c";
            when x"04b" => mem_addr <= x"09d";
            when x"00d" => mem_addr <= x"09e";
            when x"04c" => mem_addr <= x"09f";
            when x"00e" => mem_addr <= x"0a0";
            when x"04d" => mem_addr <= x"0a1";
            when x"00f" => mem_addr <= x"0a2";
            when x"04e" => mem_addr <= x"0a3";
            when x"010" => mem_addr <= x"0a4";
            when x"04f" => mem_addr <= x"0a5";
            when x"011" => mem_addr <= x"0a6";
            when x"050" => mem_addr <= x"0a7";
            when x"012" => mem_addr <= x"0a8";
            when x"051" => mem_addr <= x"0a9";
            when x"013" => mem_addr <= x"0aa";
            when x"052" => mem_addr <= x"0ab";
            when x"014" => mem_addr <= x"0ac";
            when x"053" => mem_addr <= x"0ad";
            when x"015" => mem_addr <= x"0ae";
            when x"054" => mem_addr <= x"0af";
            when x"016" => mem_addr <= x"0b0";
            when x"055" => mem_addr <= x"0b1";
            when x"017" => mem_addr <= x"0b2";
            when x"056" => mem_addr <= x"0b3";
            when x"018" => mem_addr <= x"0b4";
            when x"057" => mem_addr <= x"0b5";
            when x"019" => mem_addr <= x"0b6";
            when x"058" => mem_addr <= x"0b7";
            when x"01a" => mem_addr <= x"0b8";
            when x"059" => mem_addr <= x"0b9";
            when x"01b" => mem_addr <= x"0ba";
            when x"05a" => mem_addr <= x"0bb";
            when x"01c" => mem_addr <= x"0bc";
            when x"05b" => mem_addr <= x"0bd";
            when x"01d" => mem_addr <= x"0be";
            when x"05c" => mem_addr <= x"0bf";
            when x"01e" => mem_addr <= x"0c0";
            when x"05d" => mem_addr <= x"0c1";
            when x"01f" => mem_addr <= x"0c2";
            when x"05e" => mem_addr <= x"0c3";
            when x"020" => mem_addr <= x"0c4";
            when x"05f" => mem_addr <= x"0c5";
            when x"021" => mem_addr <= x"0c6";
            when x"060" => mem_addr <= x"0c7";
            when x"022" => mem_addr <= x"0c8";
            when x"061" => mem_addr <= x"0c9";
            when x"023" => mem_addr <= x"0ca";
            when x"062" => mem_addr <= x"0cb";
            when x"024" => mem_addr <= x"0cc";
            when x"063" => mem_addr <= x"0cd";
            when x"025" => mem_addr <= x"0ce";
            when x"064" => mem_addr <= x"0cf";
            when x"026" => mem_addr <= x"0d0";
            when x"065" => mem_addr <= x"0d1";
            when x"027" => mem_addr <= x"0d2";
            when x"066" => mem_addr <= x"0d3";
            when x"028" => mem_addr <= x"0d4";
            when x"067" => mem_addr <= x"0d5";
            when x"029" => mem_addr <= x"0d6";
            when x"068" => mem_addr <= x"0d7";
            when x"02a" => mem_addr <= x"0d8";
            when x"069" => mem_addr <= x"0d9";
            when x"02b" => mem_addr <= x"0da";
            when x"06a" => mem_addr <= x"0db";
            when x"02c" => mem_addr <= x"0dc";
            when x"06b" => mem_addr <= x"0dd";
            when x"02d" => mem_addr <= x"0de";
            when x"06c" => mem_addr <= x"0df";
            when x"02e" => mem_addr <= x"0e0";
            when x"06d" => mem_addr <= x"0e1";
            when x"02f" => mem_addr <= x"0e2";
            when x"06e" => mem_addr <= x"0e3";
            when x"030" => mem_addr <= x"0e4";
            when x"06f" => mem_addr <= x"0e5";
            when x"031" => mem_addr <= x"0e6";
            when x"070" => mem_addr <= x"0e7";
            when x"032" => mem_addr <= x"0e8";
            when x"071" => mem_addr <= x"0e9";
            when x"033" => mem_addr <= x"0ea";
            when x"072" => mem_addr <= x"0eb";
            when x"034" => mem_addr <= x"0ec";
            when x"073" => mem_addr <= x"0ed";
            when x"035" => mem_addr <= x"0ee";
            when x"074" => mem_addr <= x"0ef";
            when x"036" => mem_addr <= x"0f0";
            when x"075" => mem_addr <= x"0f1";
            when x"037" => mem_addr <= x"0f2";
            when x"076" => mem_addr <= x"0f3";
            when x"038" => mem_addr <= x"0f4";
            when x"077" => mem_addr <= x"0f5";
            when x"039" => mem_addr <= x"0f6";
            when x"078" => mem_addr <= x"0f7";
            when x"03a" => mem_addr <= x"0f8";
            when x"079" => mem_addr <= x"0f9";
            when x"03b" => mem_addr <= x"0fa";
            when x"07a" => mem_addr <= x"0fb";
            when x"03c" => mem_addr <= x"0fc";
            when x"07b" => mem_addr <= x"0fd";
            when x"03d" => mem_addr <= x"0fe";
            when x"07c" => mem_addr <= x"0ff";
            when x"171" => mem_addr <= x"100";
            when x"1b3" => mem_addr <= x"101";
            when x"172" => mem_addr <= x"102";
            when x"1b4" => mem_addr <= x"103";
            when x"173" => mem_addr <= x"104";
            when x"1b5" => mem_addr <= x"105";
            when x"174" => mem_addr <= x"106";
            when x"1b6" => mem_addr <= x"107";
            when x"175" => mem_addr <= x"108";
            when x"1b7" => mem_addr <= x"109";
            when x"176" => mem_addr <= x"10a";
            when x"1b8" => mem_addr <= x"10b";
            when x"177" => mem_addr <= x"10c";
            when x"1b9" => mem_addr <= x"10d";
            when x"178" => mem_addr <= x"10e";
            when x"1ba" => mem_addr <= x"10f";
            when x"179" => mem_addr <= x"110";
            when x"1bb" => mem_addr <= x"111";
            when x"17a" => mem_addr <= x"112";
            when x"1bc" => mem_addr <= x"113";
            when x"17b" => mem_addr <= x"114";
            when x"1bd" => mem_addr <= x"115";
            when x"17c" => mem_addr <= x"116";
            when x"1be" => mem_addr <= x"117";
            when x"17d" => mem_addr <= x"118";
            when x"1bf" => mem_addr <= x"119";
            when x"17e" => mem_addr <= x"11a";
            when x"1c0" => mem_addr <= x"11b";
            when x"17f" => mem_addr <= x"11c";
            when x"1c1" => mem_addr <= x"11d";
            when x"180" => mem_addr <= x"11e";
            when x"1c2" => mem_addr <= x"11f";
            when x"181" => mem_addr <= x"120";
            when x"1c3" => mem_addr <= x"121";
            when x"182" => mem_addr <= x"122";
            when x"1c4" => mem_addr <= x"123";
            when x"183" => mem_addr <= x"124";
            when x"1c5" => mem_addr <= x"125";
            when x"184" => mem_addr <= x"126";
            when x"1c6" => mem_addr <= x"127";
            when x"185" => mem_addr <= x"128";
            when x"1c7" => mem_addr <= x"129";
            when x"186" => mem_addr <= x"12a";
            when x"1c8" => mem_addr <= x"12b";
            when x"187" => mem_addr <= x"12c";
            when x"1c9" => mem_addr <= x"12d";
            when x"188" => mem_addr <= x"12e";
            when x"1ca" => mem_addr <= x"12f";
            when x"189" => mem_addr <= x"130";
            when x"1cb" => mem_addr <= x"131";
            when x"18a" => mem_addr <= x"132";
            when x"1cc" => mem_addr <= x"133";
            when x"18b" => mem_addr <= x"134";
            when x"1cd" => mem_addr <= x"135";
            when x"18c" => mem_addr <= x"136";
            when x"1ce" => mem_addr <= x"137";
            when x"18d" => mem_addr <= x"138";
            when x"1cf" => mem_addr <= x"139";
            when x"18e" => mem_addr <= x"13a";
            when x"1d0" => mem_addr <= x"13b";
            when x"18f" => mem_addr <= x"13c";
            when x"1d1" => mem_addr <= x"13d";
            when x"190" => mem_addr <= x"13e";
            when x"1d2" => mem_addr <= x"13f";
            when x"191" => mem_addr <= x"140";
            when x"1d3" => mem_addr <= x"141";
            when x"192" => mem_addr <= x"142";
            when x"1d4" => mem_addr <= x"143";
            when x"193" => mem_addr <= x"144";
            when x"1d5" => mem_addr <= x"145";
            when x"194" => mem_addr <= x"146";
            when x"1d6" => mem_addr <= x"147";
            when x"195" => mem_addr <= x"148";
            when x"1d7" => mem_addr <= x"149";
            when x"196" => mem_addr <= x"14a";
            when x"1d8" => mem_addr <= x"14b";
            when x"197" => mem_addr <= x"14c";
            when x"1d9" => mem_addr <= x"14d";
            when x"198" => mem_addr <= x"14e";
            when x"1da" => mem_addr <= x"14f";
            when x"199" => mem_addr <= x"150";
            when x"1db" => mem_addr <= x"151";
            when x"19a" => mem_addr <= x"152";
            when x"1dc" => mem_addr <= x"153";
            when x"19b" => mem_addr <= x"154";
            when x"1dd" => mem_addr <= x"155";
            when x"19c" => mem_addr <= x"156";
            when x"1de" => mem_addr <= x"157";
            when x"19d" => mem_addr <= x"158";
            when x"1df" => mem_addr <= x"159";
            when x"19e" => mem_addr <= x"15a";
            when x"1e0" => mem_addr <= x"15b";
            when x"19f" => mem_addr <= x"15c";
            when x"1e1" => mem_addr <= x"15d";
            when x"1a0" => mem_addr <= x"15e";
            when x"1e2" => mem_addr <= x"15f";
            when x"1a1" => mem_addr <= x"160";
            when x"1e3" => mem_addr <= x"161";
            when x"1a2" => mem_addr <= x"162";
            when x"1e4" => mem_addr <= x"163";
            when x"1a3" => mem_addr <= x"164";
            when x"1e5" => mem_addr <= x"165";
            when x"1a4" => mem_addr <= x"166";
            when x"1e6" => mem_addr <= x"167";
            when x"1a5" => mem_addr <= x"168";
            when x"1e7" => mem_addr <= x"169";
            when x"1a6" => mem_addr <= x"16a";
            when x"1e8" => mem_addr <= x"16b";
            when x"1a7" => mem_addr <= x"16c";
            when x"1e9" => mem_addr <= x"16d";
            when x"1a8" => mem_addr <= x"16e";
            when x"1ea" => mem_addr <= x"16f";
            when x"1a9" => mem_addr <= x"170";
            when x"1eb" => mem_addr <= x"171";
            when x"1aa" => mem_addr <= x"172";
            when x"1ec" => mem_addr <= x"173";
            when x"1ab" => mem_addr <= x"174";
            when x"1ed" => mem_addr <= x"175";
            when x"1ac" => mem_addr <= x"176";
            when x"1ee" => mem_addr <= x"177";
            when x"1ad" => mem_addr <= x"178";
            when x"1ef" => mem_addr <= x"179";
            when x"1ae" => mem_addr <= x"17a";
            when x"1f0" => mem_addr <= x"17b";
            when x"1af" => mem_addr <= x"17c";
            when x"1f1" => mem_addr <= x"17d";
            when x"1b0" => mem_addr <= x"17e";
            when x"1f2" => mem_addr <= x"17f";
            when x"1b1" => mem_addr <= x"180";
            when x"1f3" => mem_addr <= x"181";
            when x"1b2" => mem_addr <= x"182";
            when x"0bb" => mem_addr <= x"183";
            when x"07d" => mem_addr <= x"184";
            when x"0bc" => mem_addr <= x"185";
            when x"07e" => mem_addr <= x"186";
            when x"0bd" => mem_addr <= x"187";
            when x"07f" => mem_addr <= x"188";
            when x"0be" => mem_addr <= x"189";
            when x"080" => mem_addr <= x"18a";
            when x"0bf" => mem_addr <= x"18b";
            when x"081" => mem_addr <= x"18c";
            when x"0c0" => mem_addr <= x"18d";
            when x"082" => mem_addr <= x"18e";
            when x"0c1" => mem_addr <= x"18f";
            when x"083" => mem_addr <= x"190";
            when x"0c2" => mem_addr <= x"191";
            when x"084" => mem_addr <= x"192";
            when x"0c3" => mem_addr <= x"193";
            when x"085" => mem_addr <= x"194";
            when x"0c4" => mem_addr <= x"195";
            when x"086" => mem_addr <= x"196";
            when x"0c5" => mem_addr <= x"197";
            when x"087" => mem_addr <= x"198";
            when x"0c6" => mem_addr <= x"199";
            when x"088" => mem_addr <= x"19a";
            when x"0c7" => mem_addr <= x"19b";
            when x"089" => mem_addr <= x"19c";
            when x"0c8" => mem_addr <= x"19d";
            when x"08a" => mem_addr <= x"19e";
            when x"0c9" => mem_addr <= x"19f";
            when x"08b" => mem_addr <= x"1a0";
            when x"0ca" => mem_addr <= x"1a1";
            when x"08c" => mem_addr <= x"1a2";
            when x"0cb" => mem_addr <= x"1a3";
            when x"08d" => mem_addr <= x"1a4";
            when x"0cc" => mem_addr <= x"1a5";
            when x"08e" => mem_addr <= x"1a6";
            when x"0cd" => mem_addr <= x"1a7";
            when x"08f" => mem_addr <= x"1a8";
            when x"0ce" => mem_addr <= x"1a9";
            when x"090" => mem_addr <= x"1aa";
            when x"0cf" => mem_addr <= x"1ab";
            when x"091" => mem_addr <= x"1ac";
            when x"0d0" => mem_addr <= x"1ad";
            when x"092" => mem_addr <= x"1ae";
            when x"0d1" => mem_addr <= x"1af";
            when x"093" => mem_addr <= x"1b0";
            when x"0d2" => mem_addr <= x"1b1";
            when x"094" => mem_addr <= x"1b2";
            when x"0d3" => mem_addr <= x"1b3";
            when x"095" => mem_addr <= x"1b4";
            when x"0d4" => mem_addr <= x"1b5";
            when x"096" => mem_addr <= x"1b6";
            when x"0d5" => mem_addr <= x"1b7";
            when x"097" => mem_addr <= x"1b8";
            when x"0d6" => mem_addr <= x"1b9";
            when x"098" => mem_addr <= x"1ba";
            when x"0d7" => mem_addr <= x"1bb";
            when x"099" => mem_addr <= x"1bc";
            when x"0d8" => mem_addr <= x"1bd";
            when x"09a" => mem_addr <= x"1be";
            when x"0d9" => mem_addr <= x"1bf";
            when x"09b" => mem_addr <= x"1c0";
            when x"0da" => mem_addr <= x"1c1";
            when x"09c" => mem_addr <= x"1c2";
            when x"0db" => mem_addr <= x"1c3";
            when x"09d" => mem_addr <= x"1c4";
            when x"0dc" => mem_addr <= x"1c5";
            when x"09e" => mem_addr <= x"1c6";
            when x"0dd" => mem_addr <= x"1c7";
            when x"09f" => mem_addr <= x"1c8";
            when x"0de" => mem_addr <= x"1c9";
            when x"0a0" => mem_addr <= x"1ca";
            when x"0df" => mem_addr <= x"1cb";
            when x"0a1" => mem_addr <= x"1cc";
            when x"0e0" => mem_addr <= x"1cd";
            when x"0a2" => mem_addr <= x"1ce";
            when x"0e1" => mem_addr <= x"1cf";
            when x"0a3" => mem_addr <= x"1d0";
            when x"0e2" => mem_addr <= x"1d1";
            when x"0a4" => mem_addr <= x"1d2";
            when x"0e3" => mem_addr <= x"1d3";
            when x"0a5" => mem_addr <= x"1d4";
            when x"0e4" => mem_addr <= x"1d5";
            when x"0a6" => mem_addr <= x"1d6";
            when x"0e5" => mem_addr <= x"1d7";
            when x"0a7" => mem_addr <= x"1d8";
            when x"0e6" => mem_addr <= x"1d9";
            when x"0a8" => mem_addr <= x"1da";
            when x"0e7" => mem_addr <= x"1db";
            when x"0a9" => mem_addr <= x"1dc";
            when x"0e8" => mem_addr <= x"1dd";
            when x"0aa" => mem_addr <= x"1de";
            when x"0e9" => mem_addr <= x"1df";
            when x"0ab" => mem_addr <= x"1e0";
            when x"0ea" => mem_addr <= x"1e1";
            when x"0ac" => mem_addr <= x"1e2";
            when x"0eb" => mem_addr <= x"1e3";
            when x"0ad" => mem_addr <= x"1e4";
            when x"0ec" => mem_addr <= x"1e5";
            when x"0ae" => mem_addr <= x"1e6";
            when x"0ed" => mem_addr <= x"1e7";
            when x"0af" => mem_addr <= x"1e8";
            when x"0ee" => mem_addr <= x"1e9";
            when x"0b0" => mem_addr <= x"1ea";
            when x"0ef" => mem_addr <= x"1eb";
            when x"0b1" => mem_addr <= x"1ec";
            when x"0f0" => mem_addr <= x"1ed";
            when x"0b2" => mem_addr <= x"1ee";
            when x"0f1" => mem_addr <= x"1ef";
            when x"0b3" => mem_addr <= x"1f0";
            when x"0f2" => mem_addr <= x"1f1";
            when x"0b4" => mem_addr <= x"1f2";
            when x"0f3" => mem_addr <= x"1f3";
            when x"0b5" => mem_addr <= x"1f4";
            when x"0f4" => mem_addr <= x"1f5";
            when x"0b6" => mem_addr <= x"1f6";
            when x"0f5" => mem_addr <= x"1f7";
            when x"0b7" => mem_addr <= x"1f8";
            when x"0f6" => mem_addr <= x"1f9";
            when x"0b8" => mem_addr <= x"1fa";
            when x"0f7" => mem_addr <= x"1fb";
            when x"0b9" => mem_addr <= x"1fc";
            when x"0f8" => mem_addr <= x"1fd";
            when x"0ba" => mem_addr <= x"1fe";
            when x"0f9" => mem_addr <= x"1ff";
            when others => mem_addr <= (others => '0');
        end case;
    end process;
end RTL;
